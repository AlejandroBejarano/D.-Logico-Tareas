`timescale 1ns/1ps

 module module_decoder_tb (

 );
    
 endmodule